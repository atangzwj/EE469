module regfile (
    output logic [63:0] ReadData1,
    output logic [63:0] ReadData2,
    input  logic [63:0] WriteData,
    input  logic [4:0]  ReadRegister1,
    input  logic [4:0]  ReadRegister2,
    input  logic [4:0]  WriteRegister,
    input               RegWrite,
    input               clk,
    );

endmodule
