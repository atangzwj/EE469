module regfile (
    output [63:0] ReadData1,
    output [63:0] ReadData2,
    input  [63:0] WriteData,
    input  [4:0]  ReadRegister1,
    input  [4:0]  ReadRegister2,
    input  [4:0]  WriteRegister,
    input         RegWrite,
    input         clk,
    );






endmodule
