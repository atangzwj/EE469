module regfile (
    output logic [0:63] ReadData1,
    output logic [0:63] ReadData2,
    input  logic [0:63] WriteData,
    input  logic [0:4]  ReadRegister1,
    input  logic [0:4]  ReadRegister2,
    input  logic [0:4]  WriteRegister,
    input  logic        RegWrite,
    input  logic        clk,
    );






endmodule
