module regfile (
    output [0:63] ReadData1,
    output [0:63] ReadData2,
    input  [0:63] WriteData,
    input  [0:4]  ReadRegister1,
    input  [0:4]  ReadRegister2,
    input  [0:4]  WriteRegister,
    input         RegWrite,
    input         clk,
    );






endmodule
