`timescale 1ns/10ps

module main_control (
   output logic reg2Loc,
   output logic ALU_src,
   output logic memToReg,
   input  logic [20:0] opcode;
   );

   
endmodule
